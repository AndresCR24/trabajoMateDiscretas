��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  A 1 N ?     W      �  � 1 � ?     X      �  � 1 ?     Y      �  i1 s?     Z                  ��� 	 CLogicOut�� 	 CTerminal  �@�A               �            �8�H           ��    ��  CNAND�  (8=9              @          �  (H=I              @          �  T@iA               �            <4TL           ��    ��  CNAND3�  �H�I                          �  �X�Y                          �  �h�i                          �  �XY              @            �D�l           ��( $   ��  � �!                          �  �0�1                          �  �()              @            ��4           ��    ��  ����               �            ����     !      ��    ��  (�=�              @          �  (�=�     	         @          �  (�=�              @          �  d�y�               �            <�d�     #      ��( $   ��  ����                          �  ����                          �  ���              @            ����     (      ��    ��  ����               �            �x��     ,      ��    ��  (p=q              @          �  (�=�              @          �  (�=�              @          �  d�y�               �            <ld�     .      ��( $   ��  ����                          �  ����              @          �  ����              @          �  ���              @            ����     3      ��( $   ��  �p�q                          �  ����                          �  �xy              @            �l��     8      ��    ��  �H�I              @          �  �X�Y                          �  �PQ              @            �D�\     <      ��    ��  �� ��                �            �� ��      @      ��    ��  (� =�               @          �  (� =�               @          �  (� =�               @          �  d� y�                �            <� d�      B      ��( $   ��  ��              @          �  � �!                          �  �0�1              @          �  � !              @            ��4     G      ��( $   ��  �� ��               @          �  �� ��               @          �  �� ��                           �  �� �               @            �� ��      L      ��( $   ��  �� ��                           �  �� ��                           �  �� �               @            �� ��      Q      ��    �� 	 CRailThru�  �p��      	 d       @          �  �t��              @            �r��    V    ����    T��  ppq�       d                   �  ptq�                            lrt�    Y    ����    �� 	 CInverter�   h !}        	                   �   � !�               @            | ,�     ]      ��    ��   T !i                             D (T     `      ��    [��  �h �}        	                   �  �� ��      	         @            || ��     b      ��    [��  � h � }        	                   �  � � � �               @            � | � �     e      ��    [��  h h i }        	                   �  h � i �               @            \ | t �     h      ��    ��  �T �i                             �D �T     k      ��    ��  � T � i                             � D � T     m      ��    ��  h T i i                             ` D p T     o      ��    T��   p�       d                   �   t�                            � r�    q    ����    T��  p�       d       @          �  t�              @            r�    t    ����    T��  � p� �       d                   �  � t� �                            � r� �    w    ����    T��  � p� �       d       @          �  � t� �     
         @            � r� �    z    ����    T��  ` pa �       d       @          �  ` ta �              @            \ rd �    }    ����    T��  H pI �       d                   �  H tI �                            D rL �    �    ����    ��  CLogicIn�� 	 CLatchKey  � I  W       �   �  T 	i                             L T     �    ����     ����  � I � W       �   �  � T � i                             � L � T     �    ����     ����  0 I @ W       �   �  H T I i                             D L L T     �    ����     ����  XI hW       �   �  pT qi                             lL tT     �    ����                 ���  CWire  h@�A      ��  HY       ��  H)I      ��   (9       ��   8)9      ��  phqq       ���� 
 CCrossOver  nDtL      ��  nTt\        p0qi       ����  �d�l        ph�i      ����  �d�l      ��  �T�\      ��  �D�L      ��  �,�4      ��  ��$      ��  ��        � �q      	 ��  � X� q       ����  � D� L        � �� Y       ����  � T� \      ��  � T\      ��  T$\      ��  nTt\      ��  �T�\        � X�Y      ����  � T� \      ��  � D� L      ��  � �� �      ��  � �� �        � �� q       ����  � T\      ��  � DL          q       ����  T$\      ��  D$L      ��  $$         !q       ��  H HI q       ��  H �I I       ����  f Dl L      ��  � D� L      ��  � D� L      ��  � DL      ��  D$L      ��  nDtL      ��  �D�L        H H�I      ����  f Dl L      ��  f �l �      ��  f �l �        h Hi q       ����  nt      ��  nt$      ��  n,t4      ��  nDtL      ��  nTt\      ��  nltt      ��  n|t�      ��  n�t�      ��  n�t�      ��  n�t�      ��  n�t�      ��  n�t�      ��  nt      ��  nt$        p� q1       ����  �,�4        p0�1      ����  � ��      ��  � ��      ��  � ��      ��  � ��         �!       ����  $$      ��  nt$      ��  ��$          �!      ����  n� t�       ��  n� t�       ��  n� t�       ��  n� t�         ph q�        ��  Pq       ��  � !       ��  x���      ����  �$�      ��  �$�         �!	       ����  nt      ��  ��         		      ��  �		       ��  �)�      ����  �� ��       ��  �� ��       ��  �� ��       ��  �� ��       ��  �� ��       ��  ��      ��  ��$      ��  �,�4      ��  �D�L      ��  �T�\      ��  �l�t      ��  �|��      ��  ����      ��  ����      ��  ����      ��  ����      ��  ����        �� �      	 ��  � �     	 ��  ���      	 ��  ��)�     	 ��   �)�      ����  � �� �      ��  � �� �        � p� �       ����  � �� �      ��  � ��      ��  �$�      ��  n�t�      ��  ����        � ���      ��  H �I �       ����  f �l �      ��  � �� �      ��  � �� �      ��  � ��      ��  �$�      ��  n�t�      ��  ����        H ���      ��  ��       ��  x���      ��  ��      ��  �)�      ��   x�       ��   �)�      ��   PQ      ��  p)q      ��  � �        ����  D$L      ��  T$\      ��  l$t      ��  |$�      ��  �$�      ��  �$�         0!�       ����  n�t�      ��  ����         ���      ����  � � � �       ��  � � � �       ��  � �       ��  � � $      ��  � D� L      ��  � T� \      ��  � l� t      ��  � �� �        � � � �       ����  � ��      ��  �$�      ��  n�t�      ��  ����        � ���      ��  H � I �       ����  f �l �      ��  � �� �      ��  � �� �      ��  � ��      ��  �$�      ��  n�t�      ��  ����        H ���      ����  � � �       ��  �       ��  � $      ��  � DL      ��  � T\      ��  � lt         � �       ����  |$�      ��  n|t�      ��  �|��         ���      ��  � X� q       ����  � l� t      ��  � lt      ��  l$t      ��  nltt      ��  �l�t        � p�q      ����  � D� L        �  � Y       ����  � T� \      ��  � T\      ��  T$\      ��  nTt\      ��  �T�\        � X�Y      ��  h i I       ����  � D� L      ��  � D� L      ��  � DL      ��  D$L      ��  nDtL      ��  �D�L        h H�I      ��  x� ��       ��   !      ��  � )�       ��  � )�       ��   � �       ��  � )�       ����  $      ��  $$         � !1       ����  n,t4      ��  �,�4         0�1      ����  � � � �       ��  � � � �       ��  � �         � h � !       ����  � � $      ��  � $      ��  $$      ��  nt$      ��  ��$        �  �!      ����  � �       ��  � �       ��  �       ��  $      ��  nt      ��  ��        h �      ��  h � i        ����  �� ��         p� ��       ����  � $�       ��  � $�       ��  � $�          � !�        ����  n� t�       ��  �� ��          � ��       ����  f � l �         h � i �        ����  � � � �       ��  � � � �       ��  � � �       ��  � $�       ��  n� t�       ��  �� ��         h � ��       ����  � � �          h �        ����  � $�       ��  n� t�       ��  �� ��          � ��       ��  H p I �        ����  f � l �       ��  � � � �       ��  � � � �       ��  � � �       ��  � $�       ��  n� t�       ��  �� ��         H � ��       ��  ph �i       ��  p!q      ��  h !i       ��   h 	i       ��  � h � i       ��  � h � i       ��  H h i i       ��  H h I q        ��  � p� q      ��  ` pi q                  �                         �   �   �    �  �   �   �    �  �   �    � ! � ! # # $ $ % � % & & � ( ( ) ) * * , , . !. / / 0 0 1 1 3 <3 4 64 5 *5 6 6 8 P8 9 K9 : : < _< = X= > >  @ f@ B kB C iC D hD E E fG |G H vH I oI J J gL �L M �M N �N O O iQ �Q R �R S S j� V W W   � Y Z Z   ] ` ] ^ ^ �` ` �b k b c c � e m e f f -h o h i i �k k �m m �o o �� q r r   �t u u   � w x x   �z { {   �} ~ ~   � � � �   � � �� � �� � �� � �  �  �   � �  � Y � � � � � � � � �  � � � � � � � � � � � � � V � w � � � � � � � � � � � � � �  � � � � � � -�� � � � � q � � � � � � � �� � � � � � � � � � � � � � � � � �  � � � � =^�� �� z� p� d� \� T� M� B� 9� +� � � � � � � � � � �  � @� 7� � D� � � � � � � �  � �� �� �� �� � !hg& ! � � #� � � � � � � � � � % � �� �� �� �� �� �� {� q� e� ]� U� N� C� :� ,� � c � $ * # >O� � � � � ) ;� 
� � � � � ( 1 , 6 0 : / > � � . jk#c#[#S#L#A#8l**� *� 5 -�-�-~-w-a-Y-Q-?f 66� 6)6� 6 � 4 �<<� <	<5<� <(<� <� 3 D�DDxDbDZDR�KK'K� K� � 9 VPP4PJP&P� P� 8 V`rXX3XIX%X� X� O= �__W_2_H_$_� _� � < E @ J � � D O C S ""B l�ly�oo� o� #I r�r�r}�vv1vGvnv� v� VH |u|0|F|m|� |� ^G �|�� � N ������^ ��� �� lM ��i ��t�/�E���� �� �L �������� �� DR �����s�.������ �� ;Q � b t � �] �� r� �e � h ��z � } �              �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 